
assign PCIE_CHNL_RX_IF = PCIE_CHNL_TX_IF;
assign PCIE_CHNL_RX_LAST_IF = PCIE_CHNL_TX_LAST_IF;
assign PCIE_CHNL_RX_LEN_IF = PCIE_CHNL_TX_LEN_IF;
assign PCIE_CHNL_RX_OFF_IF = PCIE_CHNL_TX_OFF_IF;
assign PCIE_CHNL_RX_DATA_IF = PCIE_CHNL_TX_DATA_IF;
assign PCIE_CHNL_RX_DATA_VALID_IF = PCIE_CHNL_TX_DATA_VALID_IF;
assign PCIE_CHNL_TX_ACK_IF = PCIE_CHNL_RX_ACK_IF;
assign PCIE_CHNL_TX_DATA_REN_IF = PCIE_CHNL_RX_DATA_REN_IF;

assign PLD_CLK_IF = PLD_CLK;


`IOB_CLOCK(PLD_CLK,16)


